module foo1;
// 20171030a, master-001
endmodule
