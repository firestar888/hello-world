module foo1;
// 20171030a, branch "readme-edits" 003
endmodule
