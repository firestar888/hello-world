module foo1;
// 20171030a, branch "readme-edits" 001
endmodule
