module foo1;
// 20171030a
endmodule
