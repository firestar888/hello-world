module foo1;
// 20171030a, master-002
endmodule
